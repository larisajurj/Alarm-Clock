module LongShortPressesdetector_tb();
endmodule
